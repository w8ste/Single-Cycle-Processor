module datapath();

endmodule // datapath
