module controller();

endmodule // controller
